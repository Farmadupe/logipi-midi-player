--library ieee;
--use ieee.std_logic_1164.all;
--use ieee.numeric_std.all;
--use ieee.math_real.all;

--library virtual_button_lib;
--use virtual_button_lib.midi_pkg.all;
--use virtual_button_lib.constants.all;
--use virtual_button_lib.utils.all;
--use virtual_button_lib.sine_lut_pkg.all;

--entity sine_generator is
--  port(
--    ctrl    : in ctrl_t;
--    midi_no : in midi_note_t;

--    sine_read_address : out integer range 0 to sine_addr_max
--    );
--end;



--architecture rtl of sine_generator is


--  -- sine signals
--  signal sine_read_address : integer range 0 to sine_addr_max;
--  signal sine_read_out     : signed(15 downto 0);

--  -- other internals
--begin





--end;
