library ieee;
use ieee.std_logic_1164.all;

library virtual_button_lib;
use virtual_button_lib.utils.all;
use virtual_button_lib.constants.all;

entity spi_enqueue_serializer is
  port();
end;

architecture rtl of spi_enqueue_serializer is
begin
end;
