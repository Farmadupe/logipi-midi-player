package constants is
  constant clk_period : time := 20 ns;

  constant spi_word_length : integer := 8;
end;
