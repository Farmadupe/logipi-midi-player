library ieee;
use ieee.std_logic_1164.all;

library virtual_button_lib;

entity midi_ram is
  generic num_brams
end;

architecture rtl of midi_ram is
begin
end;
