package uart_constants is
  constant baud_rate : integer := 9600;
end;
