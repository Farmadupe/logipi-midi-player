package uart_constants is
  constant baud_rate : integer := 115200;
end;
